// Button/Switch Output Module
// input
// the button raw values
// output
// the fancy fancy flip flopped, filtered outputs

module input_filtering (
    input  [3:0] buttonRaw,
    output [3:0] buttonFiltered
);


endmodule  //button_output
